`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   23:13:23 10/22/2020
// Design Name:   four_one_mux
// Module Name:   /home/ise/Xilinx_Shared/Lab1/four_one_mux_test.v
// Project Name:  Lab1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: four_one_mux
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module four_one_mux_test;

	// Outputs
	//wire ;

	// Instantiate the Unit Under Test (UUT)
	/*four_one_mux uut (
		.()
	);*/

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

